
module nios_system (
	clk_clk,
	reset_reset_n,
	switches_export);	

	input		clk_clk;
	input		reset_reset_n;
	input		switches_export;
endmodule
